// 64bit floating point multiplier testbench  

`include "fp-mult.v"

module multiplier_tb ();

    reg [63:0] A, B;
    wire [63:0] out;
    
	initial begin
        A = 64'b1_10000000000_0000000000000000000000000000000000000000000000000000;//-2.00
		B = 64'b0_01111111111_0000000000000000000000000000000000000000000000000000;//1.00
        #5;

        A = 64'b1_11111111111_0000000000000000000000000000000000000000000000000000;   // infi
		B = 64'b0_01111111111_0000000000000000000000000000000000000000000000000000;//1.00
        #5;

        A = 64'b0_10000000101_0000011111101100101111111011000101011011010101110011;  // 65.9812
        B = 64'b0_10000000101_0100100001111101111100111011011001000101101000011100;  // 82.123
        // ans = 0_10000001011_0101001010101001001011110111011001111010101100001000
        #5;
        
        A = 64'b1_00000000000_0000000000000000000000000000000000000000000000000000;//-2.00
		B = 64'b0_01111111111_0000000000000000000000000000000000000000000000000000;//1.00
        #5;

        $finish;
    end

	double_multiplier d1(A, B, out);
    initial begin
        $monitor(" A = %b\n B = %b\n out = %b_%b_%b\n", A, B, out[63], out[62:52], out[51:0]);
    end
    
endmodule

