// 64bit floating point adder testbench  

`include "FPAdder.v"

module fpadder_tb();
    reg [63:0] a, b;
    wire [63:0] out;

    initial begin

        a=64'b0_11111111111_0111001100110011001100110011001100110011001100110011;			// 1.45
		b=64'b0_11111111111_1000110011001100110011001100110011001100110011001101;			// 1.55
		// ans = 0_10000000000_1000000000000000000000000000000000000000000000000000         
		#10;

        a=64'b0_01111111111_0000000000000000000000000000000000000000000000000000;			// 1.00
        b=64'b0_10000000000_0000000000000000000000000000000000000000000000000000;			// 2.00
		// ans = 0_10000000000_1000000000000000000000000000000000000000000000000000   
		#10;

		a=64'b1_10000001100_0001100001000110001111010111000010100011110101110001;	//-8968.78
		b=64'b0_10000001101_1100101010001111100000100000110001001001101110100110;	//29347.877
		// ans = 0_10000001101_0011111001101100011000110101001111110111110011101110  20379.097
		#10;

		a=64'b1_10000001100_0011000110010101010111000010100011110101110000101000;    // -9778.67
		b=64'b0_10000001100_0011000110010101010111000010100011110101110000101000;    // 9778.67
		// ans = 0 ,  0
		#10;


        // /////  this one is wrong...
		a=64'b0_01111111111_0111001100110011001100110011001100110011001100110011;			// 1.45
		b=64'b1_01111111111_1000110011001100110011001100110011001100110011001100;			// -1.55
		// ans = 1_01111111011_1001100110011001100110011001100110011001100110010000
		#10;

		a=64'b1_01111111111_0111001100110011001100110011001100110011001100110011;			// -1.45
		b=64'b1_01111111111_1000110011001100110011001100110011001100110011001100;			// -1.55
		// ans = 1_10000000000_0111111111111111111111111111111111111111111111111111
		#10;


		a=64'b0_01111111111_0000000000000000000000000000000000000000000000000000;			// 1.00
		b=64'b1_10000000000_0000000000000000000000000000000000000000000000000000;			// -2.00
		// ans = 1_01111111111_0000000000000000000000000000000000000000000000000000;
		#10;

		$finish; 

    end

    fp_adder FP1 (a, b, out);


    initial begin
        $monitor("output: %b %b %b", out[63], out[62:52], out[51:0]);
    end

endmodule


