// recursive adder testbench....

`include "adder_64.v"

module adder_tb();
    reg [63:0] a,b;
    reg cin;
    wire [63:0] sum;
	wire cout;

    initial begin
        a = 64'b000000000000000000000000000000000000000000000000000000000010101;  // 21
		b = 64'b000000000000000000000000000000000000000000000000000000000010100;  // 20
        cin = 0;
        #5;

        a = 64'b000000000000000000000000000000000000000000000000000000011000000;  // 192
		b = 64'b000000000000000000000000000000000000000000000000000000000001000;  // 8
        cin = 0;
        #5;

        a = 64'b000000000000000000000000000000000000000000000000110010001110000;  // 25712
		b = 64'b000000000000000000000000000000000000101011111101001011010010011;  // 92182163
        cin = 0;
        #5;

        a = 64'b000000000000000000000000000000000000000000000000000000000000000;  // 0
		b = 64'b000000000000000000000000000000000000101011111101001011010010011;  // 92182163
        cin = 0;
        #5;

        a = 64'b111111111111111111111111111111111111111111111111111111111111111;  // infinity
		b = 64'b000000000000000000000000000000000000101011111101001011010010011;  // 92182163
        cin = 0;
        #5;

        $finish;
    end

    adder_64bit a1(a, b, cin, sum, cout);
    initial begin
        $monitor(" a = %d b = %d cin = %b\n out = %d cout = %b\n", a, b, cin, sum, cout);
    end

endmodule


