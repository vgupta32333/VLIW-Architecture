// wallace tree multiplier test bench..
`include "WTM.v"

module wallace_tb ();
    reg [63:0] a, b;
    wire [127:0] out;

    initial begin
        a = 64'b0000000000000000000000000000000000000000000000000000000000001011;  // 11
		b = 64'b0000000000000000000000000000000000000000000000000000000000010100;  // 20
        #5;

        a = 64'b0000000000000000000000000000000000000000000000000000000000000000;  // 0
		b = 64'b0000000000000000000000000000000000000000000000000000000000010100;  // 20
        #5;

        a = 64'b1111111111111111111111111111111111111111111111111111111111111111;  
		b = 64'b1111111111111111111111111111111111111111111111111111111111111111;  
        #5;

        a = 64'b0000000000000000000000000000000000000000000000000000001101101100;  // 876
		b = 64'b0000000000000000000000000000000000000000000000000000010001000100;  // 1092
        #5;

        a = 64'b0000000000000000000000000000000000000000000011101001100010110000;  // 956592
		b = 64'b0000000000000000000000000000000000000000100010000001010011010111;  // 8918231
        #5;

        $finish;
    end

    wallace_64bit w1(a, b, out);
    initial begin
        $monitor(" a = %d\n b = %d\n out = %b", a, b, out);
    end

endmodule
